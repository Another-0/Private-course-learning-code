`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:38:00 06/16/2021 
// Design Name: 
// Module Name:    yumeng2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module yumeng2(a,b,c
    );
	 input a,b;
	 output c;
	 assign c = a&b;

endmodule
